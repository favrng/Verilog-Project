// hallo.v
module hallo;
  initial 
    begin
      $display("Hallo Sayang ...");
      $finish ;
    end
endmodule
